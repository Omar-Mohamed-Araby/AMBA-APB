module Top (PCLK,PRESETn,MADDR,MWDATA,MSTRB,MWRITE,MREQ,MPROT,MSLVERR,MRDATA,MREADY);

    parameter ADDR_WIDTH = 32;
    parameter DATA_WIDTH = 32;
    parameter STROBE_WIDTH = DATA_WIDTH/8;
    parameter PROT_WIDTH = 3;

    input PCLK,PRESETn;
    input [PROT_WIDTH-1:0] MPROT;
    input [ADDR_WIDTH-1:0] MADDR;
    input MWRITE;
    input MREQ;
    input [DATA_WIDTH-1:0] MWDATA;
    input [STROBE_WIDTH-1:0] MSTRB;


    output MSLVERR;
    output [DATA_WIDTH-1:0] MRDATA;
    output MREADY;

    wire [ADDR_WIDTH-1:0] PADDR;
    wire PSEL0,PSEL1;
    wire [PROT_WIDTH-1:0] PPROT;
    wire PWRITE;
    wire [DATA_WIDTH-1:0] PWDATA;
    wire [STROBE_WIDTH-1:0] PSTRB;
    wire PENABLE;
    wire PREADY;
    wire PSLVERR;
    wire [DATA_WIDTH-1:0] PRDATA;
    wire PREADY0,PREADY1;
    wire [DATA_WIDTH-1:0] PRDATA0,PRDATA1;
    wire PSLVERR0,PSLVERR1;
    wire LPSEL0 ,LPSEL1;

    assign PREADY  = (PSEL0) ? PREADY0  : (PSEL1) ? PREADY1  : 1'b0;

    assign PRDATA  = (LPSEL0) ? PRDATA0  : (LPSEL1) ? PRDATA1  : 'b0;

    assign PSLVERR = (LPSEL0) ? PSLVERR0 : (LPSEL1) ? PSLVERR1 : 1'b0;


    APB_BUS APB (PCLK,PRESETn,PADDR,PPROT,PSEL0,PSEL1,PENABLE,PWRITE,PWDATA,PSTRB,PREADY,PRDATA,PSLVERR,
    MADDR,MWDATA,MSTRB,MWRITE,MREQ,MPROT,MSLVERR,MRDATA,MREADY);


   SLAVE_WRAPPER slave1 (PCLK,PRESETn,PADDR,PPROT,PSEL0,PENABLE,PWRITE,PWDATA,PSTRB,PREADY0,PRDATA0,PSLVERR0,LPSEL0);

   SLAVE_WRAPPER slave2 (PCLK,PRESETn,PADDR,PPROT,PSEL1,PENABLE,PWRITE,PWDATA,PSTRB,PREADY1,PRDATA1,PSLVERR1,LPSEL1);
    
endmodule